`timescale 1ns / 1ps

module skid_buffer #(parameter DWIDTH = 8)
                    (input                   i_clock,
                     input                   i_areset_n,
                     input  [(DWIDTH - 1):0] i_data,
                     input                   i_data_valid,
                     output                  o_data_ready,
                     output [(DWIDTH - 1):0] o_data,
                     output                  o_data_valid,
                     input                   i_data_ready);

  reg [(DWIDTH - 1):0] reg_data;
  reg [(DWIDTH - 1):0] next_data;

  reg                  reg_data_ready;
  reg                  next_data_ready;

  reg                  reg_bypass;
  reg                  next_bypass;

  wire                 stall;
  wire                 hand_shake;

  always @(posedge i_clock, negedge i_areset_n)
    if (~i_areset_n)
      begin
        reg_data       <= {DWIDTH{1'b0}};
        reg_data_ready <= 1'b0;
        reg_bypass     <= 1'b1;
      end
    else
      begin
        reg_data       <= next_data;
        reg_data_ready <= next_data_ready;
        reg_bypass     <= next_bypass;
      end

  assign hand_shake = ( i_data_valid  & reg_data_ready );
  assign stall      = ( !i_data_ready & hand_shake     );

  always @(*)
    if (reg_bypass)
      begin
        next_data       = ( stall ? i_data : {DWIDTH{1'b0}} );
        next_data_ready = ( stall ? 1'b0   : 1'b1           );
        next_bypass     = ( stall ? 1'b0   : reg_bypass     );
      end
    else
      begin
        next_data       = reg_data;
        next_data_ready = ( i_data_ready ? 1'b1 : reg_data_ready );
        next_bypass     = ( i_data_ready ? 1'b1 : reg_bypass     );
      end

  assign o_data_ready = reg_data_ready;
  assign o_data_valid = ( reg_bypass ? hand_shake : 1'b1     );
  assign o_data       = ( reg_bypass ? i_data     : reg_data );

endmodule
