package axi4l_test;

  `include "test-lib/axi4l-bfm.sv"
  `include "test-lib/test-config.sv"
  `include "test-lib/transaction.sv"
  `include "test-lib/monitor.sv"
  `include "test-lib/scoreboard.sv"
  `include "test-lib/driver.sv"
  `include "test-lib/generator.sv"
  `include "test-lib/environment.sv"

endpackage
